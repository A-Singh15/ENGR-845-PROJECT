`timescale 1ns/1ps

`define SMEM_MAX 1024
`define RMEM_MAX 256
`define TRANSACTION_COUNT 10
`define DRIV_IF memoryInterface.DriverInterface.Driver_cb
`define MON_IF memoryInterface.MonitorInterface.Monitor_cb
